/*
* @file pic24_top.sv
* @brief top-level file for the PIC24
* @author Nicholas Amore namore7@gmail.com
* @date Created 12/29/2022
*/

`timescale 1ns / 100ps

module hex_sequencing_computer_top
(
	input logic i_clk_50M,
	input logic i_rstn
	
);

endmodule